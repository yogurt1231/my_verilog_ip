// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: GB_Gray_RAM_MUX.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 15.0.1 Build 150 06/03/2015 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus II License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module GB_Gray_RAM_MUX (
	data0x,
	data1x,
	sel,
	result);

	parameter	DATA_WIDTH = 30;

	input	[DATA_WIDTH-1:0]  data0x;
	input	[DATA_WIDTH-1:0]  data1x;
	input	  sel;
	output	[DATA_WIDTH-1:0]  result;

	wire [DATA_WIDTH-1:0] sub_wire5;
	wire [DATA_WIDTH-1:0] sub_wire2 = data1x[DATA_WIDTH-1:0];
	wire [DATA_WIDTH-1:0] sub_wire0 = data0x[DATA_WIDTH-1:0];
	wire [2*DATA_WIDTH-1:0] sub_wire1 = {sub_wire2, sub_wire0};
	wire  sub_wire3 = sel;
	wire  sub_wire4 = sub_wire3;
	wire [DATA_WIDTH-1:0] result = sub_wire5[DATA_WIDTH-1:0];

	lpm_mux	LPM_MUX_component (
				.data (sub_wire1),
				.sel (sub_wire4),
				.result (sub_wire5)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_size = 2,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = DATA_WIDTH,
		LPM_MUX_component.lpm_widths = 1;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "2"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "30"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
// Retrieval info: USED_PORT: data0x 0 0 30 0 INPUT NODEFVAL "data0x[29..0]"
// Retrieval info: USED_PORT: data1x 0 0 30 0 INPUT NODEFVAL "data1x[29..0]"
// Retrieval info: USED_PORT: result 0 0 30 0 OUTPUT NODEFVAL "result[29..0]"
// Retrieval info: USED_PORT: sel 0 0 0 0 INPUT NODEFVAL "sel"
// Retrieval info: CONNECT: @data 0 0 30 0 data0x 0 0 30 0
// Retrieval info: CONNECT: @data 0 0 30 30 data1x 0 0 30 0
// Retrieval info: CONNECT: @sel 0 0 1 0 sel 0 0 0 0
// Retrieval info: CONNECT: result 0 0 30 0 @result 0 0 30 0
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX.bsf TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL Gray_RAM_MUX_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
